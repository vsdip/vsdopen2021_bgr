magic
tech sky130A
timestamp 1634630016
<< nwell >>
rect 34 9234 129 9334
<< pwell >>
rect 4509 1907 4522 2009
rect 4508 1244 4521 1346
rect 4508 600 4521 702
rect 4508 6 4521 57
<< psubdiff >>
rect -589 9689 4998 9708
rect -589 9630 -349 9689
rect 4802 9630 4998 9689
rect -589 9608 4998 9630
rect -589 9504 -489 9608
rect -589 8909 -572 9504
rect -503 8909 -489 9504
rect -589 8517 -489 8909
rect -589 7922 -574 8517
rect -505 7922 -489 8517
rect -589 7483 -489 7922
rect -589 6888 -573 7483
rect -504 6888 -489 7483
rect -589 6357 -489 6888
rect -589 5762 -575 6357
rect -506 5762 -489 6357
rect -589 5278 -489 5762
rect -589 4683 -577 5278
rect -508 4683 -489 5278
rect -589 4042 -489 4683
rect -589 3447 -575 4042
rect -506 3447 -489 4042
rect -589 2461 -489 3447
rect -589 1866 -568 2461
rect -499 1866 -489 2461
rect -589 925 -489 1866
rect -589 330 -574 925
rect -505 330 -489 925
rect -589 -27 -489 330
rect 4898 9504 4998 9608
rect 4898 8909 4915 9504
rect 4984 8909 4998 9504
rect 4898 8517 4998 8909
rect 4898 7922 4913 8517
rect 4982 7922 4998 8517
rect 4898 7483 4998 7922
rect 4898 6888 4914 7483
rect 4983 6888 4998 7483
rect 4898 6357 4998 6888
rect 4898 5762 4912 6357
rect 4981 5762 4998 6357
rect 4898 5278 4998 5762
rect 4898 4683 4910 5278
rect 4979 4683 4998 5278
rect 4898 4042 4998 4683
rect 4898 3447 4912 4042
rect 4981 3447 4998 4042
rect 4898 2461 4998 3447
rect 4898 1866 4919 2461
rect 4988 1866 4998 2461
rect 4898 925 4998 1866
rect 4898 330 4913 925
rect 4982 330 4998 925
rect 4898 -27 4998 330
rect -589 -55 4998 -27
rect -589 -104 -427 -55
rect 4816 -104 4998 -55
rect -589 -127 4998 -104
<< psubdiffcont >>
rect -349 9630 4802 9689
rect -572 8909 -503 9504
rect -574 7922 -505 8517
rect -573 6888 -504 7483
rect -575 5762 -506 6357
rect -577 4683 -508 5278
rect -575 3447 -506 4042
rect -568 1866 -499 2461
rect -574 330 -505 925
rect 4915 8909 4984 9504
rect 4913 7922 4982 8517
rect 4914 6888 4983 7483
rect 4912 5762 4981 6357
rect 4910 4683 4979 5278
rect 4912 3447 4981 4042
rect 4919 1866 4988 2461
rect 4913 330 4982 925
rect -427 -104 4816 -55
<< locali >>
rect -589 9689 4998 9708
rect -589 9630 -349 9689
rect 4802 9630 4998 9689
rect -589 9608 4998 9630
rect -589 9504 -489 9608
rect -589 8909 -572 9504
rect -503 8909 -489 9504
rect -472 9565 16 9570
rect -472 9475 -467 9565
rect -367 9475 16 9565
rect 4898 9504 4998 9608
rect -472 9470 16 9475
rect 4781 9475 4915 9504
rect 34 9318 129 9334
rect 34 9249 45 9318
rect 118 9249 129 9318
rect 34 9234 129 9249
rect 4781 8954 4804 9475
rect 4857 8954 4915 9475
rect 4781 8909 4915 8954
rect 4984 8909 4998 9504
rect -589 8517 -489 8909
rect 3072 8688 3272 8698
rect 3072 8608 3082 8688
rect 3262 8608 3272 8688
rect 3072 8598 3272 8608
rect -589 7922 -574 8517
rect -505 7922 -489 8517
rect 34 8570 4010 8580
rect 34 8490 3772 8570
rect 3952 8490 4010 8570
rect 34 8480 4010 8490
rect 4898 8517 4998 8909
rect -101 8160 16 8176
rect -101 8092 -87 8160
rect -2 8092 16 8160
rect -101 8076 16 8092
rect -589 7483 -489 7922
rect -589 6888 -573 7483
rect -504 6888 -489 7483
rect -589 6357 -489 6888
rect 4898 7922 4913 8517
rect 4982 7922 4998 8517
rect 4898 7483 4998 7922
rect 4898 6888 4914 7483
rect 4983 6888 4998 7483
rect 2309 6440 2394 6722
rect 4048 6717 4881 6722
rect 4048 6627 4786 6717
rect 4876 6627 4881 6717
rect 4048 6622 4881 6627
rect -589 5762 -575 6357
rect -506 5762 -489 6357
rect 2231 6410 2308 6420
rect 2231 6328 2240 6410
rect 2301 6328 2308 6410
rect 2231 6320 2308 6328
rect 4898 6357 4998 6888
rect 4022 6154 4881 6168
rect 4022 6083 4795 6154
rect 4870 6083 4881 6154
rect 4022 6068 4881 6083
rect -589 5278 -489 5762
rect -589 4683 -577 5278
rect -508 4683 -489 5278
rect -589 4042 -489 4683
rect 4898 5762 4912 6357
rect 4981 5762 4998 6357
rect 4898 5278 4998 5762
rect 4898 4683 4910 5278
rect 4979 4683 4998 5278
rect 621 4496 728 4570
rect 1679 4569 1818 4585
rect 1679 4501 1692 4569
rect 1797 4501 1818 4569
rect 1679 4485 1818 4501
rect 603 4368 3972 4468
rect -589 3447 -575 4042
rect -506 3447 -489 4042
rect -589 2461 -489 3447
rect 4898 4042 4998 4683
rect 4898 3447 4912 4042
rect 4981 3447 4998 4042
rect 603 2875 3972 2888
rect 603 2799 3877 2875
rect 3961 2799 3972 2875
rect 603 2788 3972 2799
rect 4457 2575 4881 2582
rect 4457 2538 4791 2575
rect 4871 2538 4881 2575
rect 4457 2531 4881 2538
rect -589 1866 -568 2461
rect -499 1866 -489 2461
rect 4898 2461 4998 3447
rect 4508 2002 4881 2009
rect 4508 1914 4792 2002
rect 4872 1914 4881 2002
rect 4508 1907 4881 1914
rect -589 925 -489 1866
rect 4898 1866 4919 2461
rect 4988 1866 4998 2461
rect 4508 1339 4881 1346
rect 4508 1251 4791 1339
rect 4871 1251 4881 1339
rect 4508 1244 4881 1251
rect -589 330 -574 925
rect -505 330 -489 925
rect 4898 925 4998 1866
rect 4508 695 4881 702
rect 4508 607 4791 695
rect 4871 607 4881 695
rect 4508 600 4881 607
rect -589 -27 -489 330
rect 4898 330 4913 925
rect 4982 330 4998 925
rect 4508 50 4881 57
rect 4508 13 4791 50
rect 4871 13 4881 50
rect 4508 6 4881 13
rect 4898 -27 4998 330
rect -589 -55 4998 -27
rect -589 -104 -427 -55
rect 4816 -104 4998 -55
rect -589 -127 4998 -104
<< viali >>
rect -467 9475 -367 9565
rect 45 9367 118 9436
rect 45 9249 118 9318
rect 4804 8954 4857 9475
rect 3082 8608 3262 8688
rect 3772 8490 3952 8570
rect -87 8212 -2 8280
rect -87 8092 -2 8160
rect 4786 6627 4876 6717
rect 3791 6521 3982 6584
rect 2240 6328 2301 6410
rect 2240 6208 2301 6290
rect 4795 6083 4870 6154
rect 618 5844 684 5916
rect 1692 4501 1797 4569
rect 616 2919 723 2994
rect 3877 2799 3961 2875
rect 4791 2538 4871 2575
rect 4792 1914 4872 2002
rect 4791 1251 4871 1339
rect 4791 607 4871 695
rect 4791 13 4871 50
<< metal1 >>
rect -472 9565 -362 9588
rect -472 9475 -467 9565
rect -367 9475 -362 9565
rect -472 -7 -362 9475
rect -342 9439 -242 9588
rect -342 9367 -330 9439
rect -254 9367 -242 9439
rect -342 8281 -242 9367
rect -342 8209 -331 8281
rect -252 8209 -242 8281
rect -342 8196 -242 8209
rect -222 9325 -122 9588
rect 34 9436 129 9452
rect 34 9367 45 9436
rect 118 9367 129 9436
rect 34 9352 129 9367
rect -222 9245 -209 9325
rect -134 9245 -122 9325
rect -342 8161 -242 8176
rect -342 8089 -331 8161
rect -252 8089 -242 8161
rect -342 1737 -242 8089
rect -222 5919 -122 9245
rect 34 9318 129 9334
rect 34 9249 45 9318
rect 118 9249 129 9318
rect 34 9234 129 9249
rect 3072 8688 3272 8698
rect 3072 8608 3082 8688
rect 3262 8608 3272 8688
rect 3072 8598 3272 8608
rect 3761 8570 4009 8580
rect 3761 8490 3772 8570
rect 3952 8490 4009 8570
rect 3761 8480 4009 8490
rect 4541 8572 4641 9588
rect 4541 8488 4551 8572
rect 4633 8488 4641 8572
rect -101 8280 16 8296
rect -101 8212 -87 8280
rect -2 8212 16 8280
rect -101 8196 16 8212
rect -101 8160 16 8176
rect -101 8092 -87 8160
rect -2 8092 16 8160
rect -101 8076 16 8092
rect 3740 6584 4021 6602
rect 3740 6521 3791 6584
rect 3982 6521 4021 6584
rect 3740 6502 4021 6521
rect 4541 6584 4641 8488
rect 4541 6515 4553 6584
rect 4628 6515 4641 6584
rect 4541 6502 4641 6515
rect 4661 8690 4761 9588
rect 4661 8607 4673 8690
rect 4752 8607 4761 8690
rect 2231 6410 2308 6420
rect 2231 6328 2240 6410
rect 2301 6328 2308 6410
rect 2231 6320 2308 6328
rect 4541 6406 4641 6482
rect 4541 6330 4553 6406
rect 4632 6330 4641 6406
rect 2231 6290 2308 6300
rect 2231 6208 2240 6290
rect 2301 6208 2308 6290
rect 2231 6200 2308 6208
rect -222 5849 -206 5919
rect -141 5849 -122 5919
rect -222 5831 -122 5849
rect 603 5916 696 5931
rect 603 5844 618 5916
rect 684 5844 696 5916
rect 603 5831 696 5844
rect -342 1496 -324 1737
rect -261 1496 -242 1737
rect -342 -7 -242 1496
rect -222 2991 -122 5811
rect 1679 4569 1818 4585
rect 1679 4501 1691 4569
rect 1797 4501 1818 4569
rect 1679 4485 1818 4501
rect 4541 4569 4641 6330
rect 4661 6292 4761 8607
rect 4661 6208 4670 6292
rect 4751 6208 4761 6292
rect 4661 6068 4761 6208
rect 4781 9475 4881 9588
rect 4781 8954 4804 9475
rect 4857 8954 4881 9475
rect 4781 6717 4881 8954
rect 4781 6627 4786 6717
rect 4876 6627 4881 6717
rect 4781 6154 4881 6627
rect 4781 6083 4795 6154
rect 4870 6083 4881 6154
rect 4541 4501 4556 4569
rect 4627 4501 4641 4569
rect -222 2917 -208 2991
rect -135 2917 -122 2991
rect -222 1094 -122 2917
rect 603 2994 734 3005
rect 603 2919 616 2994
rect 723 2919 734 2994
rect 603 2905 734 2919
rect 3862 2875 3972 2888
rect 3862 2799 3877 2875
rect 3961 2799 3972 2875
rect 3862 2788 3972 2799
rect 4541 2009 4641 4501
rect 4661 2876 4761 6050
rect 4661 2801 4675 2876
rect 4750 2801 4761 2876
rect 4661 2009 4761 2801
rect 4781 2575 4881 6083
rect 4781 2538 4791 2575
rect 4871 2538 4881 2575
rect 4541 1990 4642 2009
rect 4661 1990 4762 2009
rect 4781 2002 4881 2538
rect 4781 1990 4792 2002
rect 4542 1907 4642 1990
rect 4662 1907 4762 1990
rect 4782 1914 4792 1990
rect 4872 1914 4881 2002
rect 4782 1907 4881 1914
rect 4662 1888 4761 1907
rect -222 850 -207 1094
rect -138 850 -122 1094
rect -222 -7 -122 850
rect 4541 -7 4641 1888
rect 4661 1733 4761 1888
rect 4661 1510 4680 1733
rect 4742 1510 4761 1733
rect 4661 1079 4761 1510
rect 4661 871 4683 1079
rect 4742 871 4761 1079
rect 4661 -7 4761 871
rect 4781 1339 4881 1888
rect 4781 1251 4791 1339
rect 4871 1251 4881 1339
rect 4781 695 4881 1251
rect 4781 607 4791 695
rect 4871 607 4881 695
rect 4781 50 4881 607
rect 4781 13 4791 50
rect 4871 13 4881 50
rect 4781 -7 4881 13
<< via1 >>
rect -330 9367 -254 9439
rect -331 8209 -252 8281
rect 45 9367 118 9436
rect -209 9245 -134 9325
rect -331 8089 -252 8161
rect 45 9249 118 9318
rect 3082 8608 3262 8688
rect 3772 8490 3952 8570
rect 4551 8488 4633 8572
rect -87 8212 -2 8280
rect -87 8092 -2 8160
rect 3791 6521 3982 6584
rect 4553 6515 4628 6584
rect 4673 8607 4752 8690
rect 2240 6328 2301 6410
rect 4553 6330 4632 6406
rect 2240 6208 2301 6290
rect -206 5849 -141 5919
rect 618 5844 684 5916
rect -324 1496 -261 1737
rect 1691 4501 1692 4569
rect 1692 4501 1797 4569
rect 4670 6208 4751 6292
rect 4556 4501 4627 4569
rect -208 2917 -135 2991
rect 616 2919 723 2994
rect 3877 2799 3961 2875
rect 4675 2801 4750 2876
rect 3444 1518 3641 1715
rect -207 850 -138 1094
rect 3444 874 3641 1071
rect 4680 1510 4742 1733
rect 4683 871 4742 1079
<< metal2 >>
rect -342 9439 129 9452
rect -342 9367 -330 9439
rect -254 9436 129 9439
rect -254 9367 45 9436
rect 118 9367 129 9436
rect -342 9352 129 9367
rect -222 9325 129 9334
rect -222 9245 -209 9325
rect -134 9318 129 9325
rect -134 9249 45 9318
rect 118 9249 129 9318
rect -134 9245 129 9249
rect -222 9234 129 9245
rect 3072 8690 4761 8698
rect 3072 8688 4673 8690
rect 3072 8608 3082 8688
rect 3262 8608 4673 8688
rect 3072 8607 4673 8608
rect 4752 8607 4761 8690
rect 3072 8598 4761 8607
rect 3761 8572 4641 8580
rect 3761 8570 4551 8572
rect 3761 8490 3772 8570
rect 3952 8490 4551 8570
rect 3761 8488 4551 8490
rect 4633 8488 4641 8572
rect 3761 8480 4641 8488
rect -342 8281 16 8296
rect -342 8209 -331 8281
rect -252 8280 16 8281
rect -252 8212 -87 8280
rect -2 8212 16 8280
rect -252 8209 16 8212
rect -342 8196 16 8209
rect -342 8161 16 8176
rect -342 8089 -331 8161
rect -252 8160 16 8161
rect -252 8092 -87 8160
rect -2 8092 16 8160
rect -252 8089 16 8092
rect -342 8076 16 8089
rect 3740 6584 4641 6602
rect 3740 6521 3791 6584
rect 3982 6521 4553 6584
rect 3740 6515 4553 6521
rect 4628 6515 4641 6584
rect 3740 6502 4641 6515
rect 2231 6410 4641 6420
rect 2231 6328 2240 6410
rect 2301 6406 4641 6410
rect 2301 6330 4553 6406
rect 4632 6330 4641 6406
rect 2301 6328 4641 6330
rect 2231 6320 4641 6328
rect 2231 6292 4761 6300
rect 2231 6290 4670 6292
rect 2231 6208 2240 6290
rect 2301 6208 4670 6290
rect 4751 6208 4761 6292
rect 2231 6200 4761 6208
rect -222 5919 696 5931
rect -222 5849 -206 5919
rect -141 5916 696 5919
rect -141 5849 618 5916
rect -222 5844 618 5849
rect 684 5844 696 5916
rect -222 5831 696 5844
rect 1679 4569 4641 4585
rect 1679 4501 1691 4569
rect 1797 4501 4556 4569
rect 4627 4501 4641 4569
rect 1679 4485 4641 4501
rect -222 2994 734 3005
rect -222 2991 616 2994
rect -222 2917 -208 2991
rect -135 2919 616 2991
rect 723 2919 734 2994
rect -135 2917 734 2919
rect -222 2905 734 2917
rect 3862 2876 4761 2888
rect 3862 2875 4675 2876
rect 3862 2799 3877 2875
rect 3961 2801 4675 2875
rect 4750 2801 4761 2876
rect 3961 2799 4761 2801
rect 3862 2788 4761 2799
rect -342 1737 2111 1760
rect -342 1496 -324 1737
rect -261 1496 2111 1737
rect -342 1473 2111 1496
rect 3399 1733 4761 1760
rect 3399 1715 4680 1733
rect 3399 1518 3444 1715
rect 3641 1518 4680 1715
rect 3399 1510 4680 1518
rect 4742 1510 4761 1733
rect 3399 1473 4761 1510
rect -222 1094 2111 1116
rect -222 850 -207 1094
rect -138 850 2111 1094
rect -222 829 2111 850
rect 3399 1079 4761 1116
rect 3399 1071 4683 1079
rect 3399 874 3444 1071
rect 3641 874 4683 1071
rect 3399 871 4683 874
rect 4742 871 4761 1079
rect 3399 829 4761 871
use pfets  pfets_0
timestamp 1634628445
transform 1 0 34 0 1 8698
box -136 -354 4112 890
use resbank  resbank_0
timestamp 1634556819
transform 1 0 599 0 1 4602
box -150 -1934 3523 1566
use pnp10  pnp10_0
timestamp 1634562067
transform 1 0 636 0 1 1282
box -649 -1289 3885 1313
use starternfet  starternfet_0
timestamp 1634207820
transform 1 0 2531 0 1 6356
box -137 -120 1626 366
use nfets  nfets_0
timestamp 1634540517
transform 1 0 309 0 1 7380
box -411 -1180 2000 916
<< labels >>
rlabel metal1 -425 9588 -425 9588 5 vdd
port 1 s
rlabel metal1 -174 9586 -174 9586 5 vref
port 2 s
rlabel metal1 -296 9582 -296 9582 1 net1
rlabel metal1 -300 8047 -300 8047 1 qp1
rlabel metal1 4832 9576 4832 9576 1 gnd
port 3 n
rlabel metal1 4698 8730 4698 8730 1 net2
rlabel metal1 -177 5791 -177 5791 1 qp3
rlabel metal1 4590 6465 4590 6465 1 rp1
rlabel metal1 4586 8749 4586 8749 1 net6
rlabel metal1 4710 2901 4710 2901 1 qp2
rlabel metal1 -435 9588 -435 9588 5 vdd
port 1 s
<< end >>
