magic
tech sky130A
timestamp 1634628445
<< nwell >>
rect -136 -354 4112 890
<< pdiff >>
rect 481 509 505 518
rect 481 28 484 509
rect 502 28 505 509
rect 481 18 505 28
rect 941 509 965 518
rect 941 28 944 509
rect 962 28 965 509
rect 941 18 965 28
rect 1861 509 1885 518
rect 1861 28 1864 509
rect 1882 28 1885 509
rect 1861 18 1885 28
rect 2321 509 2345 518
rect 2321 28 2324 509
rect 2342 28 2345 509
rect 2321 18 2345 28
rect 2551 509 2575 518
rect 2551 28 2554 509
rect 2572 28 2575 509
rect 2551 18 2575 28
rect 2781 509 2805 518
rect 2781 28 2784 509
rect 2802 28 2805 509
rect 2781 18 2805 28
rect 3241 509 3265 518
rect 3241 28 3244 509
rect 3262 28 3265 509
rect 3241 18 3265 28
rect 3471 509 3495 518
rect 3471 28 3474 509
rect 3492 28 3495 509
rect 3471 18 3495 28
rect 3931 509 3955 518
rect 3931 28 3934 509
rect 3952 28 3955 509
rect 3931 18 3955 28
<< pdiffc >>
rect 484 28 502 509
rect 944 28 962 509
rect 1864 28 1882 509
rect 2324 28 2342 509
rect 2554 28 2572 509
rect 2784 28 2802 509
rect 3244 28 3262 509
rect 3474 28 3492 509
rect 3934 28 3952 509
<< nsubdiff >>
rect -118 864 4094 872
rect -118 782 -8 864
rect 3986 782 4094 864
rect -118 772 4094 782
rect -118 762 -18 772
rect -118 -228 -109 762
rect -28 -228 -18 762
rect 3994 763 4094 772
rect -118 -236 -18 -228
rect 3994 -227 4004 763
rect 4085 -227 4094 763
rect 3994 -236 4094 -227
rect -118 -245 4094 -236
rect -118 -327 -10 -245
rect 3984 -327 4094 -245
rect -118 -336 4094 -327
<< nsubdiffcont >>
rect -8 782 3986 864
rect -109 -228 -28 762
rect 4004 -227 4085 763
rect -10 -327 3984 -245
<< poly >>
rect 48 -10 248 5
rect 48 -90 58 -10
rect 238 -90 248 -10
rect 48 -100 248 -90
rect 278 -10 478 5
rect 278 -90 288 -10
rect 468 -90 478 -10
rect 278 -100 478 -90
rect 508 -10 708 5
rect 508 -90 518 -10
rect 698 -90 708 -10
rect 508 -100 708 -90
rect 738 -10 938 5
rect 738 -90 748 -10
rect 928 -90 938 -10
rect 738 -100 938 -90
rect 968 -10 1168 5
rect 968 -90 978 -10
rect 1158 -90 1168 -10
rect 968 -100 1168 -90
rect 1198 -10 1398 5
rect 1198 -90 1208 -10
rect 1388 -90 1398 -10
rect 1198 -100 1398 -90
rect 1428 -10 1628 5
rect 1428 -90 1438 -10
rect 1618 -90 1628 -10
rect 1428 -100 1628 -90
rect 1658 -10 1858 5
rect 1658 -90 1668 -10
rect 1848 -90 1858 -10
rect 1658 -100 1858 -90
rect 1888 -10 2088 5
rect 1888 -90 1898 -10
rect 2078 -90 2088 -10
rect 1888 -100 2088 -90
rect 2118 -10 2318 5
rect 2118 -90 2128 -10
rect 2308 -90 2318 -10
rect 2118 -100 2318 -90
rect 2348 -10 2548 5
rect 2348 -90 2358 -10
rect 2538 -90 2548 -10
rect 2348 -100 2548 -90
rect 2578 -10 2778 5
rect 2578 -90 2588 -10
rect 2768 -90 2778 -10
rect 2578 -100 2778 -90
rect 2808 -10 3008 5
rect 2808 -90 2818 -10
rect 2998 -90 3008 -10
rect 2808 -100 3008 -90
rect 3038 -10 3238 5
rect 3038 -90 3048 -10
rect 3228 -90 3238 -10
rect 3038 -100 3238 -90
rect 3268 -10 3468 5
rect 3268 -90 3278 -10
rect 3458 -90 3468 -10
rect 3268 -100 3468 -90
rect 3498 -128 3698 5
rect 3498 -208 3508 -128
rect 3688 -208 3698 -128
rect 3498 -218 3698 -208
rect 3728 -128 3928 5
rect 3728 -208 3738 -128
rect 3918 -208 3928 -128
rect 3728 -218 3928 -208
<< polycont >>
rect 58 -90 238 -10
rect 288 -90 468 -10
rect 518 -90 698 -10
rect 748 -90 928 -10
rect 978 -90 1158 -10
rect 1208 -90 1388 -10
rect 1438 -90 1618 -10
rect 1668 -90 1848 -10
rect 1898 -90 2078 -10
rect 2128 -90 2308 -10
rect 2358 -90 2538 -10
rect 2588 -90 2768 -10
rect 2818 -90 2998 -10
rect 3048 -90 3228 -10
rect 3278 -90 3458 -10
rect 3508 -208 3688 -128
rect 3738 -208 3918 -128
<< locali >>
rect -118 864 4094 872
rect -118 782 -8 864
rect 3986 782 4094 864
rect -118 772 4094 782
rect -118 762 -18 772
rect -118 -228 -109 762
rect -28 -228 -18 762
rect 3994 763 4094 772
rect 0 745 3976 754
rect 0 744 3474 745
rect 0 664 1174 744
rect 1192 664 2554 744
rect 2572 665 3474 744
rect 3492 744 3976 745
rect 3492 665 3934 744
rect 2572 664 3934 665
rect 3952 664 3976 744
rect 0 654 3976 664
rect 0 536 3976 636
rect 714 518 732 536
rect 3014 518 3032 536
rect 484 509 502 518
rect 484 18 502 28
rect 944 509 962 518
rect 1864 509 1882 518
rect 944 18 962 28
rect 1864 18 1882 28
rect 2324 509 2342 518
rect 2324 18 2342 28
rect 2554 509 2572 518
rect 2554 18 2572 28
rect 2784 509 2802 518
rect 2784 18 2802 28
rect 3244 509 3262 518
rect 3244 18 3262 28
rect 3474 509 3492 518
rect 3474 18 3492 28
rect 3934 509 3952 518
rect 3934 18 3952 28
rect 1634 0 1652 18
rect 2094 0 2112 18
rect 3704 0 3722 18
rect 3994 0 4004 763
rect 0 -10 3238 0
rect 0 -90 58 -10
rect 238 -90 288 -10
rect 468 -90 518 -10
rect 698 -90 748 -10
rect 928 -90 978 -10
rect 1158 -90 1208 -10
rect 1388 -90 1438 -10
rect 1618 -90 1668 -10
rect 1848 -90 1898 -10
rect 2078 -90 2128 -10
rect 2308 -90 2358 -10
rect 2538 -90 2588 -10
rect 2768 -90 2818 -10
rect 2998 -90 3048 -10
rect 3228 -90 3238 -10
rect 0 -100 3238 -90
rect 3268 -10 4004 0
rect 3268 -90 3278 -10
rect 3458 -90 4004 -10
rect 3268 -100 4004 -90
rect 0 -128 3976 -118
rect 0 -208 24 -128
rect 42 -208 3508 -128
rect 3688 -208 3738 -128
rect 3918 -208 3976 -128
rect 0 -218 3976 -208
rect -118 -236 -18 -228
rect 3994 -227 4004 -100
rect 4085 -227 4094 763
rect 3994 -236 4094 -227
rect -118 -245 4094 -236
rect -118 -327 -10 -245
rect 3984 -327 4094 -245
rect -118 -336 4094 -327
<< viali >>
rect 484 782 502 862
rect 944 782 962 862
rect 1404 782 1422 862
rect 1864 782 1882 862
rect 2324 782 2342 862
rect 2784 782 2802 862
rect 3244 782 3262 862
rect 1174 664 1192 744
rect 2554 664 2572 744
rect 3474 665 3492 745
rect 3934 664 3952 744
rect 24 28 42 509
rect 484 28 502 509
rect 944 28 962 509
rect 1174 28 1192 509
rect 1404 28 1422 509
rect 1864 28 1882 509
rect 2324 28 2342 509
rect 2554 28 2572 509
rect 2784 28 2802 509
rect 3244 28 3262 509
rect 3474 28 3492 509
rect 3934 28 3952 509
rect 24 -208 42 -128
<< metal1 >>
rect 481 862 505 872
rect 481 782 484 862
rect 502 782 505 862
rect 21 509 45 518
rect 21 28 24 509
rect 42 28 45 509
rect 21 -128 45 28
rect 481 509 505 782
rect 481 28 484 509
rect 502 28 505 509
rect 481 18 505 28
rect 941 862 965 872
rect 941 782 944 862
rect 962 782 965 862
rect 941 509 965 782
rect 1401 862 1425 872
rect 1401 782 1404 862
rect 1422 782 1425 862
rect 941 28 944 509
rect 962 28 965 509
rect 941 18 965 28
rect 1171 744 1195 754
rect 1171 664 1174 744
rect 1192 664 1195 744
rect 1171 509 1195 664
rect 1171 28 1174 509
rect 1192 28 1195 509
rect 1171 18 1195 28
rect 1401 509 1425 782
rect 1401 28 1404 509
rect 1422 28 1425 509
rect 1401 18 1425 28
rect 1861 862 1885 872
rect 1861 782 1864 862
rect 1882 782 1885 862
rect 1861 509 1885 782
rect 1861 28 1864 509
rect 1882 28 1885 509
rect 1861 18 1885 28
rect 2321 862 2345 872
rect 2321 782 2324 862
rect 2342 782 2345 862
rect 2321 509 2345 782
rect 2781 862 2805 872
rect 2781 782 2784 862
rect 2802 782 2805 862
rect 2321 28 2324 509
rect 2342 28 2345 509
rect 2321 18 2345 28
rect 2551 744 2575 754
rect 2551 664 2554 744
rect 2572 664 2575 744
rect 2551 509 2575 664
rect 2551 28 2554 509
rect 2572 28 2575 509
rect 2551 18 2575 28
rect 2781 509 2805 782
rect 2781 28 2784 509
rect 2802 28 2805 509
rect 2781 18 2805 28
rect 3241 862 3265 872
rect 3241 782 3244 862
rect 3262 782 3265 862
rect 3241 509 3265 782
rect 3241 28 3244 509
rect 3262 28 3265 509
rect 3241 18 3265 28
rect 3471 745 3495 754
rect 3471 665 3474 745
rect 3492 665 3495 745
rect 3471 509 3495 665
rect 3471 28 3474 509
rect 3492 28 3495 509
rect 3471 18 3495 28
rect 3931 744 3955 754
rect 3931 664 3934 744
rect 3952 664 3955 744
rect 3931 509 3955 664
rect 3931 28 3934 509
rect 3952 28 3955 509
rect 3931 18 3955 28
rect 21 -208 24 -128
rect 42 -208 45 -128
rect 21 -218 45 -208
use pfet  pfet_1
timestamp 1634550790
transform 1 0 278 0 1 18
box -48 -18 248 518
use pfet  pfet_0
timestamp 1634550790
transform 1 0 48 0 1 18
box -48 -18 248 518
use pfet  pfet_2
timestamp 1634550790
transform 1 0 508 0 1 18
box -48 -18 248 518
use pfet  pfet_3
timestamp 1634550790
transform 1 0 738 0 1 18
box -48 -18 248 518
use pfet  pfet_5
timestamp 1634550790
transform 1 0 1198 0 1 18
box -48 -18 248 518
use pfet  pfet_4
timestamp 1634550790
transform 1 0 968 0 1 18
box -48 -18 248 518
use pfet  pfet_6
timestamp 1634550790
transform 1 0 1428 0 1 18
box -48 -18 248 518
use pfet  pfet_7
timestamp 1634550790
transform 1 0 1658 0 1 18
box -48 -18 248 518
use pfet  pfet_8
timestamp 1634550790
transform 1 0 1888 0 1 18
box -48 -18 248 518
use pfet  pfet_9
timestamp 1634550790
transform 1 0 2118 0 1 18
box -48 -18 248 518
use pfet  pfet_10
timestamp 1634550790
transform 1 0 2348 0 1 18
box -48 -18 248 518
use pfet  pfet_11
timestamp 1634550790
transform 1 0 2578 0 1 18
box -48 -18 248 518
use pfet  pfet_12
timestamp 1634550790
transform 1 0 2808 0 1 18
box -48 -18 248 518
use pfet  pfet_14
timestamp 1634550790
transform 1 0 3268 0 1 18
box -48 -18 248 518
use pfet  pfet_13
timestamp 1634550790
transform 1 0 3038 0 1 18
box -48 -18 248 518
use pfet  pfet_15
timestamp 1634550790
transform 1 0 3498 0 1 18
box -48 -18 248 518
use pfet  pfet_16
timestamp 1634550790
transform 1 0 3728 0 1 18
box -48 -18 248 518
<< labels >>
rlabel locali 8 -51 8 -51 1 net2
port 4 n
rlabel locali 19 707 19 707 1 net1
port 2 n
rlabel locali 25 586 25 586 1 vref
port 3 n
rlabel locali 7 -151 7 -151 1 net6
port 5 n
rlabel locali -64 825 -64 825 1 vdd
port 6 n
<< end >>
