magic
tech sky130A
timestamp 1634207820
<< psubdiff >>
rect -137 357 1626 366
rect -137 276 -18 357
rect 1509 276 1626 357
rect -137 266 1626 276
rect -137 257 -28 266
rect -137 -10 -129 257
rect -38 -10 -28 257
rect 1517 257 1626 266
rect -137 -20 -28 -10
rect 1517 -10 1527 257
rect 1618 -10 1626 257
rect 1517 -20 1626 -10
rect -137 -30 1626 -20
rect -137 -111 -18 -30
rect 1509 -111 1626 -30
rect -137 -120 1626 -111
<< psubdiffcont >>
rect -18 276 1509 357
rect -129 -10 -38 257
rect 1527 -10 1618 257
rect -18 -111 1509 -30
<< poly >>
rect 44 236 716 246
rect 44 156 54 236
rect 706 156 716 236
rect 44 126 716 156
rect 774 236 1446 246
rect 774 156 784 236
rect 1436 156 1446 236
rect 774 126 1446 156
<< polycont >>
rect 54 156 706 236
rect 784 156 1436 236
<< locali >>
rect -137 357 1626 366
rect -137 276 -18 357
rect 1509 276 1626 357
rect -137 266 1626 276
rect -137 257 -28 266
rect -137 -10 -129 257
rect -38 113 -28 257
rect 1517 257 1626 266
rect 0 236 754 246
rect 0 156 54 236
rect 706 156 754 236
rect 0 146 754 156
rect 774 236 1490 246
rect 774 156 784 236
rect 1436 156 1490 236
rect 774 146 1490 156
rect 736 113 754 146
rect 1466 113 1484 146
rect -38 13 6 113
rect -38 -10 -28 13
rect -137 -20 -28 -10
rect 1517 -10 1527 257
rect 1618 -10 1626 257
rect 1517 -20 1626 -10
rect -137 -30 1626 -20
rect -137 -111 -18 -30
rect 1509 -111 1626 -30
rect -137 -120 1626 -111
use nfet1  nfet1_1
timestamp 1634205135
transform 1 0 760 0 1 13
box -30 -13 730 113
use nfet1  nfet1_0
timestamp 1634205135
transform 1 0 30 0 1 13
box -30 -13 730 113
<< labels >>
rlabel locali 1474 199 1474 199 1 net6
port 1 n
rlabel locali -121 328 -121 328 1 gnd
port 2 n
<< end >>
