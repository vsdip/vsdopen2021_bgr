magic
tech sky130A
timestamp 1634556819
<< pwell >>
rect -150 -1934 3523 1566
<< psubdiff >>
rect -150 1556 3523 1566
rect -150 1476 4 1556
rect 3373 1476 3523 1556
rect -150 1466 3523 1476
rect -150 1212 -50 1466
rect 3423 1212 3523 1466
rect -150 -1580 -141 1212
rect -60 -1580 -50 1212
rect -150 -1834 -50 -1580
rect 3423 -1580 3433 1212
rect 3514 -1580 3523 1212
rect 3423 -1834 3523 -1580
rect -150 -1844 3523 -1834
rect -150 -1924 4 -1844
rect 3373 -1924 3523 -1844
rect -150 -1934 3523 -1924
<< psubdiffcont >>
rect 4 1476 3373 1556
rect -141 -1580 -60 1212
rect 3433 -1580 3514 1212
rect 4 -1924 3373 -1844
<< xpolycontact >>
rect 2156 996 2297 1212
rect 814 10 949 206
rect 1083 -574 1218 -376
rect 1083 -1570 1218 -1372
<< locali >>
rect -150 1556 3523 1566
rect -150 1476 4 1556
rect 3373 1476 3523 1556
rect -150 1466 3523 1476
rect -150 1212 -50 1466
rect 4 1436 3373 1446
rect 4 1356 1083 1436
rect 1218 1356 2159 1436
rect 2294 1356 3373 1436
rect 4 1346 3373 1356
rect 4 1229 683 1329
rect 811 1319 1490 1329
rect 811 1239 814 1319
rect 949 1239 1490 1319
rect 811 1229 1490 1239
rect -150 -1580 -141 1212
rect -60 996 145 1212
rect 273 996 414 1229
rect 1349 1212 1490 1229
rect 1618 1229 2424 1329
rect 2552 1319 3373 1329
rect 2552 1239 3107 1319
rect 3229 1239 3373 1319
rect 2552 1229 3373 1239
rect 542 996 811 1212
rect 1618 996 1759 1229
rect 1887 996 2028 1229
rect 2425 996 2835 1212
rect 2963 996 3104 1229
rect 3423 1212 3523 1466
rect 3232 996 3433 1212
rect -60 216 -50 996
rect 3423 216 3433 996
rect -60 0 145 216
rect 273 0 683 216
rect 811 206 952 216
rect 811 10 814 206
rect 949 10 952 206
rect 811 0 952 10
rect 1349 0 1759 216
rect 2694 0 3104 216
rect 3373 0 3433 216
rect -60 -368 -50 0
rect 1080 -17 1221 0
rect 1887 -17 2028 0
rect 2425 -17 2566 0
rect 4 -117 1221 -17
rect 1348 -117 3364 -17
rect 4 -144 3373 -134
rect 4 -224 1083 -144
rect 1218 -224 2159 -144
rect 2294 -224 3373 -144
rect 4 -234 3373 -224
rect 4 -351 2425 -251
rect 2566 -261 3373 -251
rect 2566 -341 3107 -261
rect 3229 -341 3373 -261
rect 2566 -351 3373 -341
rect 811 -368 952 -351
rect 1349 -368 1490 -351
rect 2963 -368 3104 -351
rect 3423 -368 3433 0
rect -60 -584 4 -368
rect 273 -584 683 -368
rect 1618 -584 2028 -368
rect 2425 -584 2835 -368
rect 3373 -584 3433 -368
rect -60 -1364 -50 -584
rect 3423 -1364 3433 -584
rect -60 -1580 4 -1364
rect 414 -1580 952 -1364
rect 1349 -1580 1759 -1364
rect 2835 -1580 2963 -1364
rect 3373 -1580 3433 -1364
rect 3514 -1580 3523 1212
rect -150 -1834 -50 -1580
rect 273 -1597 414 -1580
rect 1887 -1597 2028 -1580
rect 2425 -1597 2566 -1580
rect 4 -1697 414 -1597
rect 542 -1697 3373 -1597
rect 4 -1724 3373 -1714
rect 4 -1804 1083 -1724
rect 1218 -1804 2159 -1724
rect 2294 -1804 3373 -1724
rect 4 -1814 3373 -1804
rect 3423 -1834 3523 -1580
rect -150 -1844 3523 -1834
rect -150 -1924 4 -1844
rect 3373 -1924 3523 -1844
rect -150 -1934 3523 -1924
<< viali >>
rect 1083 1356 1218 1436
rect 2159 1356 2294 1436
rect 814 1239 949 1319
rect 3107 1239 3229 1319
rect 1083 1006 1218 1202
rect 2159 1006 2294 1202
rect 814 10 949 206
rect 2159 10 2294 206
rect 1083 -224 1218 -144
rect 2159 -224 2294 -144
rect 3107 -341 3229 -261
rect 1083 -574 1218 -376
rect 2159 -576 2294 -378
rect 1083 -1570 1218 -1372
rect 2159 -1570 2294 -1374
rect 1083 -1804 1218 -1724
rect 2159 -1804 2294 -1724
<< metal1 >>
rect 1080 1436 1221 1446
rect 1080 1356 1083 1436
rect 1218 1356 1221 1436
rect 811 1319 952 1329
rect 811 1239 814 1319
rect 949 1239 952 1319
rect 811 206 952 1239
rect 1080 1202 1221 1356
rect 1080 1006 1083 1202
rect 1218 1006 1221 1202
rect 1080 996 1221 1006
rect 2156 1436 2297 1446
rect 2156 1356 2159 1436
rect 2294 1356 2297 1436
rect 2156 1202 2297 1356
rect 2156 1006 2159 1202
rect 2294 1006 2297 1202
rect 2156 996 2297 1006
rect 3104 1319 3232 1329
rect 3104 1239 3107 1319
rect 3229 1239 3232 1319
rect 811 10 814 206
rect 949 10 952 206
rect 811 0 952 10
rect 2156 206 2297 216
rect 2156 10 2159 206
rect 2294 10 2297 206
rect 1080 -144 1221 -134
rect 1080 -224 1083 -144
rect 1218 -224 1221 -144
rect 1080 -376 1221 -224
rect 1080 -574 1083 -376
rect 1218 -574 1221 -376
rect 1080 -584 1221 -574
rect 2156 -144 2297 10
rect 2156 -224 2159 -144
rect 2294 -224 2297 -144
rect 2156 -378 2297 -224
rect 3104 -261 3232 1239
rect 3104 -341 3107 -261
rect 3229 -341 3232 -261
rect 3104 -351 3232 -341
rect 2156 -576 2159 -378
rect 2294 -576 2297 -378
rect 2156 -584 2297 -576
rect 1080 -1372 1221 -1364
rect 1080 -1570 1083 -1372
rect 1218 -1570 1221 -1372
rect 1080 -1724 1221 -1570
rect 1080 -1804 1083 -1724
rect 1218 -1804 1221 -1724
rect 1080 -1814 1221 -1804
rect 2156 -1374 2297 -1364
rect 2156 -1570 2159 -1374
rect 2294 -1570 2297 -1374
rect 2156 -1724 2297 -1570
rect 2156 -1804 2159 -1724
rect 2294 -1804 2297 -1724
rect 2156 -1814 2297 -1804
use res1p41  res1p41_13
timestamp 1633868552
transform 1 0 4 0 1 -1364
box -4 -216 145 996
use res1p41  res1p41_14
timestamp 1633868552
transform 1 0 273 0 1 -1364
box -4 -216 145 996
use res1p41  res1p41_16
timestamp 1633868552
transform 1 0 811 0 1 -1364
box -4 -216 145 996
use res1p41  res1p41_15
timestamp 1633868552
transform 1 0 542 0 1 -1364
box -4 -216 145 996
use res1p41  res1p41_17
timestamp 1633868552
transform 1 0 1080 0 1 -1364
box -4 -216 145 996
use res1p41  res1p41_19
timestamp 1633868552
transform 1 0 1618 0 1 -1364
box -4 -216 145 996
use res1p41  res1p41_18
timestamp 1633868552
transform 1 0 1349 0 1 -1364
box -4 -216 145 996
use res1p41  res1p41_20
timestamp 1633868552
transform 1 0 1887 0 1 -1364
box -4 -216 145 996
use res1p41  res1p41_22
timestamp 1633868552
transform 1 0 2425 0 1 -1364
box -4 -216 145 996
use res1p41  res1p41_21
timestamp 1633868552
transform 1 0 2156 0 1 -1364
box -4 -216 145 996
use res1p41  res1p41_23
timestamp 1633868552
transform 1 0 2694 0 1 -1364
box -4 -216 145 996
use res1p41  res1p41_25
timestamp 1633868552
transform 1 0 3232 0 1 -1364
box -4 -216 145 996
use res1p41  res1p41_24
timestamp 1633868552
transform 1 0 2963 0 1 -1364
box -4 -216 145 996
use res1p41  res1p41_0
timestamp 1633868552
transform 1 0 4 0 1 216
box -4 -216 145 996
use res1p41  res1p41_1
timestamp 1633868552
transform 1 0 273 0 1 216
box -4 -216 145 996
use res1p41  res1p41_2
timestamp 1633868552
transform 1 0 542 0 1 216
box -4 -216 145 996
use res1p41  res1p41_3
timestamp 1633868552
transform 1 0 811 0 1 216
box -4 -216 145 996
use res1p41  res1p41_4
timestamp 1633868552
transform 1 0 1080 0 1 216
box -4 -216 145 996
use res1p41  res1p41_5
timestamp 1633868552
transform 1 0 1349 0 1 216
box -4 -216 145 996
use res1p41  res1p41_6
timestamp 1633868552
transform 1 0 1618 0 1 216
box -4 -216 145 996
use res1p41  res1p41_7
timestamp 1633868552
transform 1 0 1887 0 1 216
box -4 -216 145 996
use res1p41  res1p41_8
timestamp 1633868552
transform 1 0 2156 0 1 216
box -4 -216 145 996
use res1p41  res1p41_9
timestamp 1633868552
transform 1 0 2425 0 1 216
box -4 -216 145 996
use res1p41  res1p41_10
timestamp 1633868552
transform 1 0 2694 0 1 216
box -4 -216 145 996
use res1p41  res1p41_11
timestamp 1633868552
transform 1 0 2963 0 1 216
box -4 -216 145 996
use res1p41  res1p41_12
timestamp 1633868552
transform 1 0 3232 0 1 216
box -4 -216 145 996
<< labels >>
rlabel locali -93 1509 -93 1509 1 gnd
port 1 n
rlabel locali 30 1284 30 1284 1 vref
port 2 n
rlabel locali 39 -1770 39 -1770 1 qp2
port 4 n
rlabel locali 47 -1652 47 -1652 1 qp3
port 5 n
rlabel locali 35 -65 35 -65 1 rp1
port 6 n
<< end >>
