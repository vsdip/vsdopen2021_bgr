magic
tech sky130A
timestamp 1634540517
<< ndiff >>
rect 263 503 287 513
rect 263 23 266 503
rect 284 23 287 503
rect 263 13 287 23
rect 1303 503 1327 513
rect 1303 23 1306 503
rect 1324 23 1327 503
rect 1303 13 1327 23
rect 1433 503 1457 513
rect 1433 23 1436 503
rect 1454 23 1457 503
rect 1433 13 1457 23
rect 1563 503 1587 513
rect 1563 23 1566 503
rect 1584 23 1587 503
rect 1563 13 1587 23
rect 1820 503 1850 513
rect 1820 23 1826 503
rect 1844 23 1850 503
rect 1820 13 1850 23
rect 263 -287 287 -277
rect 263 -767 266 -287
rect 284 -767 287 -287
rect 263 -777 287 -767
rect 1303 -287 1327 -277
rect 1303 -767 1306 -287
rect 1324 -767 1327 -287
rect 1303 -777 1327 -767
rect 1433 -287 1457 -277
rect 1433 -767 1436 -287
rect 1454 -767 1457 -287
rect 1433 -777 1457 -767
rect 1563 -287 1587 -277
rect 1563 -767 1566 -287
rect 1584 -767 1587 -287
rect 1563 -777 1587 -767
<< ndiffc >>
rect 266 23 284 503
rect 1306 23 1324 503
rect 1436 23 1454 503
rect 1566 23 1584 503
rect 1826 23 1844 503
rect 266 -767 284 -287
rect 1306 -767 1324 -287
rect 1436 -767 1454 -287
rect 1566 -767 1584 -287
<< psubdiff >>
rect -410 666 2000 676
rect -410 586 -300 666
rect 1890 586 2000 666
rect -410 576 2000 586
rect -410 566 -310 576
rect -410 -830 -400 566
rect -320 -830 -310 566
rect 1900 566 2000 576
rect -410 -840 -310 -830
rect 1900 -830 1910 566
rect 1990 -830 2000 566
rect 1900 -840 2000 -830
rect -410 -850 2000 -840
rect -410 -930 -300 -850
rect 1890 -930 2000 -850
rect -410 -940 2000 -930
<< psubdiffcont >>
rect -300 586 1890 666
rect -400 -830 -320 566
rect 1910 -830 1990 566
rect -300 -930 1890 -850
<< poly >>
rect -230 -25 -130 0
rect -230 -55 -220 -25
rect -140 -55 -130 -25
rect -230 -209 -130 -55
rect -230 -239 -220 -209
rect -140 -239 -130 -209
rect -230 -264 -130 -239
rect -100 -25 0 0
rect -100 -55 -91 -25
rect -11 -55 0 -25
rect -100 -209 0 -55
rect -100 -239 -90 -209
rect -10 -239 0 -209
rect -100 -264 0 -239
rect 30 -92 130 0
rect 30 -172 40 -92
rect 120 -172 130 -92
rect 30 -264 130 -172
rect 160 -92 260 0
rect 160 -172 170 -92
rect 250 -172 260 -92
rect 160 -264 260 -172
rect 290 -25 390 0
rect 290 -55 300 -25
rect 380 -55 390 -25
rect 290 -209 390 -55
rect 290 -239 300 -209
rect 380 -239 390 -209
rect 290 -264 390 -239
rect 420 -25 520 0
rect 420 -55 430 -25
rect 509 -55 520 -25
rect 420 -209 520 -55
rect 420 -239 430 -209
rect 509 -239 520 -209
rect 420 -264 520 -239
rect 550 -92 650 0
rect 550 -172 560 -92
rect 640 -172 650 -92
rect 550 -264 650 -172
rect 680 -92 780 0
rect 680 -172 690 -92
rect 770 -172 780 -92
rect 680 -264 780 -172
rect 810 -92 910 0
rect 810 -172 820 -92
rect 900 -172 910 -92
rect 810 -264 910 -172
rect 940 -92 1040 0
rect 940 -172 950 -92
rect 1030 -172 1040 -92
rect 940 -264 1040 -172
rect 1070 -25 1170 0
rect 1070 -55 1081 -25
rect 1160 -55 1170 -25
rect 1070 -209 1170 -55
rect 1070 -239 1081 -209
rect 1160 -239 1170 -209
rect 1070 -264 1170 -239
rect 1200 -25 1300 0
rect 1200 -55 1210 -25
rect 1290 -55 1300 -25
rect 1200 -209 1300 -55
rect 1200 -239 1210 -209
rect 1290 -239 1300 -209
rect 1200 -264 1300 -239
rect 1330 -92 1430 0
rect 1330 -172 1340 -92
rect 1420 -172 1430 -92
rect 1330 -264 1430 -172
rect 1460 -92 1560 0
rect 1460 -172 1470 -92
rect 1550 -172 1560 -92
rect 1460 -264 1560 -172
rect 1590 -25 1690 0
rect 1590 -55 1600 -25
rect 1680 -55 1690 -25
rect 1590 -209 1690 -55
rect 1590 -239 1601 -209
rect 1681 -239 1690 -209
rect 1590 -264 1690 -239
rect 1720 -25 1820 0
rect 1720 -55 1730 -25
rect 1810 -55 1820 -25
rect 1720 -209 1820 -55
rect 1720 -239 1730 -209
rect 1810 -239 1820 -209
rect 1720 -264 1820 -239
<< polycont >>
rect -220 -55 -140 -25
rect -220 -239 -140 -209
rect -91 -55 -11 -25
rect -90 -239 -10 -209
rect 40 -172 120 -92
rect 170 -172 250 -92
rect 300 -55 380 -25
rect 300 -239 380 -209
rect 430 -55 509 -25
rect 430 -239 509 -209
rect 560 -172 640 -92
rect 690 -172 770 -92
rect 820 -172 900 -92
rect 950 -172 1030 -92
rect 1081 -55 1160 -25
rect 1081 -239 1160 -209
rect 1210 -55 1290 -25
rect 1210 -239 1290 -209
rect 1340 -172 1420 -92
rect 1470 -172 1550 -92
rect 1600 -55 1680 -25
rect 1601 -239 1681 -209
rect 1730 -55 1810 -25
rect 1730 -239 1810 -209
<< locali >>
rect -410 906 2000 916
rect -410 826 -257 906
rect -233 826 136 906
rect 154 905 1436 906
rect 154 826 717 905
rect 735 826 1436 905
rect 1454 826 1823 906
rect 1847 826 2000 906
rect -410 816 2000 826
rect -410 786 2000 796
rect -410 706 6 786
rect 24 706 266 786
rect 284 706 916 786
rect 934 706 1306 786
rect 1324 706 1566 786
rect 1584 706 2000 786
rect -410 696 2000 706
rect -410 666 2000 676
rect -410 586 -300 666
rect 1890 586 2000 666
rect -410 576 2000 586
rect -410 566 -310 576
rect -410 -830 -400 566
rect -320 -15 -310 566
rect -254 513 -236 576
rect -124 513 -106 576
rect 396 513 414 576
rect 656 551 934 556
rect 656 534 851 551
rect 868 534 934 551
rect 656 532 934 534
rect 656 513 674 532
rect 916 513 934 532
rect 1176 513 1194 576
rect 1696 513 1714 576
rect 266 503 284 513
rect 266 13 284 23
rect 1306 503 1324 513
rect 1306 13 1324 23
rect 1436 503 1454 513
rect 1436 13 1454 23
rect 1566 503 1584 513
rect 1566 13 1584 23
rect 1826 503 1844 576
rect 1826 13 1844 23
rect 1900 566 2000 576
rect 526 -15 544 13
rect 786 -15 804 13
rect 1046 -15 1064 13
rect 1900 -15 1910 566
rect -320 -25 509 -15
rect -320 -55 -220 -25
rect -140 -55 -91 -25
rect -11 -55 300 -25
rect 380 -55 430 -25
rect -320 -65 509 -55
rect 526 -24 1064 -15
rect 526 -56 656 -24
rect 674 -56 1064 -24
rect 526 -65 1064 -56
rect 1081 -25 1910 -15
rect 1160 -55 1210 -25
rect 1290 -55 1600 -25
rect 1680 -55 1730 -25
rect 1810 -55 1910 -25
rect 1081 -65 1910 -55
rect -320 -199 -310 -65
rect -260 -92 1850 -82
rect -260 -172 -257 -92
rect -233 -172 40 -92
rect 120 -172 170 -92
rect 250 -172 560 -92
rect 640 -172 690 -92
rect 770 -172 820 -92
rect 900 -172 950 -92
rect 1030 -172 1340 -92
rect 1420 -172 1470 -92
rect 1550 -172 1823 -92
rect 1847 -172 1850 -92
rect -260 -182 1850 -172
rect 1900 -199 1910 -65
rect -320 -209 509 -199
rect -320 -239 -220 -209
rect -140 -239 -90 -209
rect -10 -239 300 -209
rect 380 -239 430 -209
rect -320 -249 509 -239
rect 526 -209 1064 -199
rect 526 -239 916 -209
rect 934 -239 1064 -209
rect 526 -249 1064 -239
rect 1081 -209 1910 -199
rect 1160 -239 1210 -209
rect 1290 -239 1601 -209
rect 1681 -239 1730 -209
rect 1810 -239 1910 -209
rect 1081 -249 1910 -239
rect -320 -830 -310 -249
rect 526 -277 544 -249
rect 786 -277 804 -249
rect 1046 -277 1064 -249
rect 266 -287 284 -277
rect 266 -777 284 -767
rect 1306 -287 1324 -277
rect 1306 -777 1324 -767
rect 1436 -287 1454 -277
rect 1436 -777 1454 -767
rect 1566 -287 1584 -277
rect 1566 -777 1584 -767
rect -410 -840 -310 -830
rect -254 -840 -236 -777
rect -124 -840 -106 -777
rect 396 -840 414 -777
rect 656 -796 674 -777
rect 916 -796 934 -777
rect 656 -798 934 -796
rect 656 -815 718 -798
rect 735 -815 934 -798
rect 656 -820 934 -815
rect 1176 -840 1194 -777
rect 1696 -840 1714 -777
rect 1826 -840 1844 -777
rect 1900 -830 1910 -249
rect 1990 -830 2000 566
rect 1900 -840 2000 -830
rect -410 -850 2000 -840
rect -410 -930 -300 -850
rect 1890 -930 2000 -850
rect -410 -940 2000 -930
rect -410 -968 2000 -960
rect -410 -1050 6 -968
rect 24 -1050 266 -968
rect 284 -969 1306 -968
rect 284 -1050 656 -969
rect -410 -1051 656 -1050
rect 674 -1050 1306 -969
rect 1324 -1050 1566 -968
rect 1584 -1050 2000 -968
rect 674 -1051 2000 -1050
rect -410 -1060 2000 -1051
rect -411 -1088 1999 -1080
rect -411 -1170 136 -1088
rect 154 -1091 1436 -1088
rect 154 -1170 850 -1091
rect 868 -1170 1436 -1091
rect 1454 -1170 1999 -1088
rect -411 -1180 1999 -1170
<< viali >>
rect -257 826 -233 906
rect 136 826 154 906
rect 717 826 735 905
rect 1436 826 1454 906
rect 1823 826 1847 906
rect 6 706 24 786
rect 266 706 284 786
rect 916 706 934 786
rect 1306 706 1324 786
rect 1566 706 1584 786
rect 851 534 868 551
rect 6 23 24 503
rect 136 23 154 503
rect 266 23 284 503
rect 1306 23 1324 503
rect 1436 23 1454 503
rect 1566 23 1584 503
rect 656 -56 674 -24
rect -257 -172 -233 -92
rect 1823 -172 1847 -92
rect 916 -239 934 -209
rect 6 -767 24 -287
rect 136 -767 154 -287
rect 266 -767 284 -287
rect 1306 -767 1324 -287
rect 1436 -767 1454 -287
rect 1566 -767 1584 -287
rect 718 -815 735 -798
rect 6 -1050 24 -968
rect 266 -1050 284 -968
rect 656 -1051 674 -969
rect 1306 -1050 1324 -968
rect 1566 -1050 1584 -968
rect 136 -1170 154 -1088
rect 850 -1170 868 -1091
rect 1436 -1170 1454 -1088
<< metal1 >>
rect -260 906 -230 916
rect -260 826 -257 906
rect -233 826 -230 906
rect -260 -92 -230 826
rect 133 906 157 916
rect 133 826 136 906
rect 154 826 157 906
rect 3 786 27 796
rect 3 706 6 786
rect 24 706 27 786
rect 3 503 27 706
rect 3 23 6 503
rect 24 23 27 503
rect 3 13 27 23
rect 133 503 157 826
rect 712 905 741 916
rect 712 826 717 905
rect 735 826 741 905
rect 133 23 136 503
rect 154 23 157 503
rect 133 13 157 23
rect 263 786 287 796
rect 263 706 266 786
rect 284 706 287 786
rect 263 503 287 706
rect 263 23 266 503
rect 284 23 287 503
rect 263 13 287 23
rect -260 -172 -257 -92
rect -233 -172 -230 -92
rect -260 -182 -230 -172
rect 653 -24 677 -15
rect 653 -56 656 -24
rect 674 -56 677 -24
rect 3 -287 27 -277
rect 3 -767 6 -287
rect 24 -767 27 -287
rect 3 -968 27 -767
rect 3 -1050 6 -968
rect 24 -1050 27 -968
rect 3 -1060 27 -1050
rect 133 -287 157 -277
rect 133 -767 136 -287
rect 154 -767 157 -287
rect 133 -1088 157 -767
rect 263 -287 287 -277
rect 263 -767 266 -287
rect 284 -767 287 -287
rect 263 -968 287 -767
rect 263 -1050 266 -968
rect 284 -1050 287 -968
rect 263 -1060 287 -1050
rect 653 -969 677 -56
rect 712 -798 741 826
rect 1433 906 1457 916
rect 1433 826 1436 906
rect 1454 826 1457 906
rect 913 786 937 796
rect 913 706 916 786
rect 934 706 937 786
rect 712 -815 718 -798
rect 735 -815 741 -798
rect 712 -820 741 -815
rect 845 551 874 556
rect 845 534 851 551
rect 868 534 874 551
rect 653 -1051 656 -969
rect 674 -1051 677 -969
rect 653 -1060 677 -1051
rect 133 -1170 136 -1088
rect 154 -1170 157 -1088
rect 133 -1180 157 -1170
rect 845 -1091 874 534
rect 913 -209 937 706
rect 1303 786 1327 796
rect 1303 706 1306 786
rect 1324 706 1327 786
rect 1303 503 1327 706
rect 1303 23 1306 503
rect 1324 23 1327 503
rect 1303 13 1327 23
rect 1433 503 1457 826
rect 1820 906 1850 916
rect 1820 826 1823 906
rect 1847 826 1850 906
rect 1433 23 1436 503
rect 1454 23 1457 503
rect 1433 13 1457 23
rect 1563 786 1587 796
rect 1563 706 1566 786
rect 1584 706 1587 786
rect 1563 503 1587 706
rect 1563 23 1566 503
rect 1584 23 1587 503
rect 1563 13 1587 23
rect 1820 -92 1850 826
rect 1820 -172 1823 -92
rect 1847 -172 1850 -92
rect 1820 -182 1850 -172
rect 913 -239 916 -209
rect 934 -239 937 -209
rect 913 -249 937 -239
rect 1303 -287 1327 -277
rect 1303 -767 1306 -287
rect 1324 -767 1327 -287
rect 1303 -968 1327 -767
rect 1303 -1050 1306 -968
rect 1324 -1050 1327 -968
rect 1303 -1060 1327 -1050
rect 1433 -287 1457 -277
rect 1433 -767 1436 -287
rect 1454 -767 1457 -287
rect 845 -1170 850 -1091
rect 868 -1170 874 -1091
rect 845 -1180 874 -1170
rect 1433 -1088 1457 -767
rect 1563 -287 1587 -277
rect 1563 -767 1566 -287
rect 1584 -767 1587 -287
rect 1563 -968 1587 -767
rect 1563 -1050 1566 -968
rect 1584 -1050 1587 -968
rect 1563 -1060 1587 -1050
rect 1433 -1170 1436 -1088
rect 1454 -1170 1457 -1088
rect 1433 -1180 1457 -1170
use nfet  nfet_31
timestamp 1634540125
transform 1 0 -230 0 1 -777
box -30 -13 130 513
use nfet  nfet_30
timestamp 1634540125
transform 1 0 -100 0 1 -777
box -30 -13 130 513
use nfet  nfet_9
timestamp 1634540125
transform 1 0 160 0 1 -777
box -30 -13 130 513
use nfet  nfet_8
timestamp 1634540125
transform 1 0 30 0 1 -777
box -30 -13 130 513
use nfet  nfet_10
timestamp 1634540125
transform 1 0 290 0 1 -777
box -30 -13 130 513
use nfet  nfet_11
timestamp 1634540125
transform 1 0 420 0 1 -777
box -30 -13 130 513
use nfet  nfet_12
timestamp 1634540125
transform 1 0 550 0 1 -777
box -30 -13 130 513
use nfet  nfet_14
timestamp 1634540125
transform 1 0 810 0 1 -777
box -30 -13 130 513
use nfet  nfet_13
timestamp 1634540125
transform 1 0 680 0 1 -777
box -30 -13 130 513
use nfet  nfet_15
timestamp 1634540125
transform 1 0 940 0 1 -777
box -30 -13 130 513
use nfet  nfet_21
timestamp 1634540125
transform 1 0 1200 0 1 -777
box -30 -13 130 513
use nfet  nfet_20
timestamp 1634540125
transform 1 0 1070 0 1 -777
box -30 -13 130 513
use nfet  nfet_22
timestamp 1634540125
transform 1 0 1330 0 1 -777
box -30 -13 130 513
use nfet  nfet_23
timestamp 1634540125
transform 1 0 1460 0 1 -777
box -30 -13 130 513
use nfet  nfet_26
timestamp 1634540125
transform 1 0 1590 0 1 -777
box -30 -13 130 513
use nfet  nfet_27
timestamp 1634540125
transform 1 0 1720 0 1 -777
box -30 -13 130 513
use nfet  nfet_29
timestamp 1634540125
transform 1 0 -230 0 1 13
box -30 -13 130 513
use nfet  nfet_28
timestamp 1634540125
transform 1 0 -100 0 1 13
box -30 -13 130 513
use nfet  nfet_0
timestamp 1634540125
transform 1 0 30 0 1 13
box -30 -13 130 513
use nfet  nfet_1
timestamp 1634540125
transform 1 0 160 0 1 13
box -30 -13 130 513
use nfet  nfet_2
timestamp 1634540125
transform 1 0 290 0 1 13
box -30 -13 130 513
use nfet  nfet_3
timestamp 1634540125
transform 1 0 420 0 1 13
box -30 -13 130 513
use nfet  nfet_4
timestamp 1634540125
transform 1 0 550 0 1 13
box -30 -13 130 513
use nfet  nfet_5
timestamp 1634540125
transform 1 0 680 0 1 13
box -30 -13 130 513
use nfet  nfet_6
timestamp 1634540125
transform 1 0 810 0 1 13
box -30 -13 130 513
use nfet  nfet_7
timestamp 1634540125
transform 1 0 940 0 1 13
box -30 -13 130 513
use nfet  nfet_17
timestamp 1634540125
transform 1 0 1200 0 1 13
box -30 -13 130 513
use nfet  nfet_16
timestamp 1634540125
transform 1 0 1070 0 1 13
box -30 -13 130 513
use nfet  nfet_18
timestamp 1634540125
transform 1 0 1330 0 1 13
box -30 -13 130 513
use nfet  nfet_19
timestamp 1634540125
transform 1 0 1460 0 1 13
box -30 -13 130 513
use nfet  nfet_24
timestamp 1634540125
transform 1 0 1590 0 1 13
box -30 -13 130 513
use nfet  nfet_25
timestamp 1634540125
transform 1 0 1720 0 1 13
box -30 -13 130 513
<< labels >>
rlabel locali -387 876 -387 876 1 net1
port 1 n
rlabel locali -378 743 -378 743 1 qp1
port 2 n
rlabel locali -367 -892 -367 -892 1 gnd
port 3 n
rlabel locali -367 -1023 -367 -1023 1 rp1
port 4 n
rlabel locali -374 -1129 -374 -1129 1 net2
port 5 n
<< end >>
